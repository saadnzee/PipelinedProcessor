module ROM_PP(
 output reg [31:0] Instr,
 input [31:0] PC_In
);

reg [31:0] memory [31:0];

initial begin 
//	WITHOUT HAZARDS
memory[0] = 32'b000000_00001_00010_10000_00000_100000; // add
memory[1] = 32'b000000_00011_00100_10001_00000_100010; // sub
memory[2] = 32'b000000_00001_00010_10011_00000_100011; // mult
memory[3] = 32'b000000_00001_00010_10011_00000_100110; // slt
memory[4] = 32'b001010_00001_00010_00000_00000_000110; // addi
memory[5] = 32'b100011_00111_10100_00000_00000_000010; // LW 
memory[6] = 32'b101011_00111_10000_00000_00000_000100; // SW 
memory[7] = 32'b000100_01000_01001_00000_00000_000110; // Branch = 6 + PC + 1 = 6+7+1 = 14
//	dummy instructions
memory[8] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[9] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[10] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[11] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[12] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[13] = 32'b000000_10000_00011_10011_00000_100000; // add
//	WITH HAZARDS (AFTER BRANCH WE COME HERE)
memory[14] = 32'b000000_00001_00011_10110_00000_100000; // add
memory[15] = 32'b000000_10110_00100_10101_00000_100010; // sub
memory[16] = 32'b000000_10110_01000_10011_00000_100100; // mult
memory[17] = 32'b100011_00111_11100_00000_00000_000011; // LW 
memory[18] = 32'b000000_11100_00011_10000_00000_100000; // add
memory[19] = 32'b100011_00110_00001_00000_00000_000010; // LW
memory[20] = 32'b100011_00001_00010_00000_00000_000010; // LW  
memory[21] = 32'b101011_00010_00111_00000_00000_000011; // SW 
memory[22] = 32'b000010_00000_00000_00000_00000_011100; // Jump
memory[23] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[24] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[25] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[26] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[27] = 32'b000000_10000_00011_10011_00000_100000; // add
memory[28] = 32'b000000_10000_00011_10011_00000_100000; // add
end

always@(*) begin
Instr <= memory[PC_In];
end

endmodule

