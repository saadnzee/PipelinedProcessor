module ROM_PP(
 output reg [31:0] Instr,
 input [31:0] PC_In
);

reg [31:0] memory [31:0];

initial begin 
// R-Type
//memory[0] = 32'b000100_01000_01001_00000_00000_001010; // Branch = 10+PC+1 = 11
memory[0] = 32'b000000_00001_00010_10000_00000_100000; // add
memory[1] = 32'b000000_10000_00100_10001_00000_100010; // sub
memory[2] = 32'b000000_10000_01000_10011_00000_100100; // mult
memory[3] = 32'b100011_00111_10100_00000_00000_000010; // LW 
//memory[4] = 32'b100011_10100_00010_00000_00000_000011; // LW
memory[4] = 32'b000000_10100_00010_10000_00000_100000; // add
// I-Type
//memory[4] = 32'b001000_00000_00001_00011_00000_100101; // addi
memory[5] = 32'b100011_00111_00100_00000_00000_000010; // LW // addr = 7, value = 5 :: rd/rt/destination = 4/100 
memory[6] = 32'b000000_00100_00001_00011_00000_100000; // R-Type ADD
memory[7] = 32'b101011_00111_00100_00000_00000_000011; // SW // add = 7, value = 5 :: 5 + 3, 8. Location 8 value saved
memory[8] = 32'b100011_00111_00101_00000_00000_000011; // LW from SW location
memory[9] = 32'b000000_00101_00001_00011_00000_100000; // R-Type ADD
memory[10] = 32'b000100_01000_01001_00000_00000_000011; // Branch = 3 + PC + 1 = 11 + 3 = 15 but instr would be 14th
memory[11] = 32'b000000_00000_00001_00100_00000_100000; // add 
memory[12] = 32'b000010_00000_00000_00000_00000_010011; // Jump
memory[13] = 32'b000000_00000_00001_00100_00000_100000; // add
memory[14] = 32'b000000_01000_00001_00101_00000_100010; // sub 
memory[15] = 32'b000000_00000_00001_00100_00000_100000; // add
memory[16] = 32'b000000_00000_00001_00100_00000_100000; // add
memory[17] = 32'b000000_00000_00001_00100_00000_100000; // add
memory[18] = 32'b000000_00000_00001_00100_00000_100000; // add
memory[19] = 32'b000000_01000_00001_00101_00000_100000; // add 
memory[20] = 32'b000000_00000_00001_00100_00000_100010; // sub (R-Type) after jump
end

always@(*) begin
Instr <= memory[PC_In];
end

endmodule

